library ieee;
use ieee.numeric_std.all;
use ieee.std_logic_1164.all;

-- Este componente es donde se almacenan las constantes de atan(2**-i) 
-- Su tama�o depende del numero de bits
-- ai -> atan(2**-i) en binario con formato punto fijo Q0.31

entity rom_atan32 is
	port(
	a0,a1,a2,a3,a4,a5,a6,a7,a8,a9,a10,a11,a12,a13,a14,a15,a16,a17,a18,a19,a20,a21,a22,a23,a24,a25,a26,a27,a28,a29,a30,a31: out signed (31 downto 0));
end entity;

architecture rtl of rom_atan32 is
type localidades is array (0 to 31) of signed (31 downto 0);
signal a: localidades:=(
"01100100100001111110110101010001",
"00111011010110001100111000001010",
"00011111010110110111010111111001",
"00001111111010101101110101001101",
"00000111111111010101011011101101",
"00000011111111111010101010110111",
"00000001111111111111010101010101",
"00000000111111111111111010101010",
"00000000011111111111111111010101",
"00000000001111111111111111111010",
"00000000000111111111111111111111",
"00000000000011111111111111111111",
"00000000000001111111111111111111",
"00000000000000111111111111111111",
"00000000000000011111111111111111",
"00000000000000001111111111111111",
"00000000000000000111111111111111",
"00000000000000000011111111111111",
"00000000000000000001111111111111",
"00000000000000000000111111111111",
"00000000000000000000011111111111",
"00000000000000000000001111111111",
"00000000000000000000000111111111",
"00000000000000000000000011111111",
"00000000000000000000000001111111",
"00000000000000000000000000111111",
"00000000000000000000000000011111",
"00000000000000000000000000010000",
"00000000000000000000000000001000",
"00000000000000000000000000000100",
"00000000000000000000000000000010",
"00000000000000000000000000000001");
begin
	a0 <= a(0);
	a1 <= a(1);
	a2 <= a(2);
	a3 <= a(3);
	a4 <= a(4);
	a5 <= a(5);
	a6 <= a(6);
	a7 <= a(7);
	a8 <= a(8);
	a9 <= a(9);
	a10 <= a(10);
	a11 <= a(11);
	a12 <= a(12);
	a13 <= a(13);
	a14 <= a(14);
	a15 <= a(15);
	a16 <= a(16);
	a17 <= a(17);
	a18 <= a(18);
	a19 <= a(19);
	a20 <= a(20);
	a21 <= a(21);
	a22 <= a(22);
	a23 <= a(23);
	a24 <= a(24);
	a25 <= a(25);
	a26 <= a(26);
	a27 <= a(27);
	a28 <= a(28);
	a29 <= a(29);
	a30 <= a(30);
	a31 <= a(31);
end rtl;